magic
tech sky130A
magscale 1 2
timestamp 1654447720
<< obsli1 >>
rect 1104 2159 68816 77809
<< obsm1 >>
rect 1104 1776 68876 77840
<< metal2 >>
rect 1306 79200 1362 80000
rect 3882 79200 3938 80000
rect 6458 79200 6514 80000
rect 9034 79200 9090 80000
rect 11610 79200 11666 80000
rect 14186 79200 14242 80000
rect 16854 79200 16910 80000
rect 19430 79200 19486 80000
rect 22006 79200 22062 80000
rect 24582 79200 24638 80000
rect 27158 79200 27214 80000
rect 29826 79200 29882 80000
rect 32402 79200 32458 80000
rect 34978 79200 35034 80000
rect 37554 79200 37610 80000
rect 40130 79200 40186 80000
rect 42706 79200 42762 80000
rect 45374 79200 45430 80000
rect 47950 79200 48006 80000
rect 50526 79200 50582 80000
rect 53102 79200 53158 80000
rect 55678 79200 55734 80000
rect 58346 79200 58402 80000
rect 60922 79200 60978 80000
rect 63498 79200 63554 80000
rect 66074 79200 66130 80000
rect 68650 79200 68706 80000
rect 1398 0 1454 800
rect 4158 0 4214 800
rect 6918 0 6974 800
rect 9770 0 9826 800
rect 12530 0 12586 800
rect 15382 0 15438 800
rect 18142 0 18198 800
rect 20994 0 21050 800
rect 23754 0 23810 800
rect 26514 0 26570 800
rect 29366 0 29422 800
rect 32126 0 32182 800
rect 34978 0 35034 800
rect 37738 0 37794 800
rect 40590 0 40646 800
rect 43350 0 43406 800
rect 46202 0 46258 800
rect 48962 0 49018 800
rect 51722 0 51778 800
rect 54574 0 54630 800
rect 57334 0 57390 800
rect 60186 0 60242 800
rect 62946 0 63002 800
rect 65798 0 65854 800
rect 68558 0 68614 800
<< obsm2 >>
rect 1418 79144 3826 79200
rect 3994 79144 6402 79200
rect 6570 79144 8978 79200
rect 9146 79144 11554 79200
rect 11722 79144 14130 79200
rect 14298 79144 16798 79200
rect 16966 79144 19374 79200
rect 19542 79144 21950 79200
rect 22118 79144 24526 79200
rect 24694 79144 27102 79200
rect 27270 79144 29770 79200
rect 29938 79144 32346 79200
rect 32514 79144 34922 79200
rect 35090 79144 37498 79200
rect 37666 79144 40074 79200
rect 40242 79144 42650 79200
rect 42818 79144 45318 79200
rect 45486 79144 47894 79200
rect 48062 79144 50470 79200
rect 50638 79144 53046 79200
rect 53214 79144 55622 79200
rect 55790 79144 58290 79200
rect 58458 79144 60866 79200
rect 61034 79144 63442 79200
rect 63610 79144 66018 79200
rect 66186 79144 68594 79200
rect 1308 856 68704 79144
rect 1308 800 1342 856
rect 1510 800 4102 856
rect 4270 800 6862 856
rect 7030 800 9714 856
rect 9882 800 12474 856
rect 12642 800 15326 856
rect 15494 800 18086 856
rect 18254 800 20938 856
rect 21106 800 23698 856
rect 23866 800 26458 856
rect 26626 800 29310 856
rect 29478 800 32070 856
rect 32238 800 34922 856
rect 35090 800 37682 856
rect 37850 800 40534 856
rect 40702 800 43294 856
rect 43462 800 46146 856
rect 46314 800 48906 856
rect 49074 800 51666 856
rect 51834 800 54518 856
rect 54686 800 57278 856
rect 57446 800 60130 856
rect 60298 800 62890 856
rect 63058 800 65742 856
rect 65910 800 68502 856
rect 68670 800 68704 856
<< metal3 >>
rect 0 78480 800 78600
rect 69200 78344 70000 78464
rect 0 75760 800 75880
rect 69200 75352 70000 75472
rect 0 73176 800 73296
rect 69200 72360 70000 72480
rect 0 70456 800 70576
rect 69200 69368 70000 69488
rect 0 67872 800 67992
rect 69200 66512 70000 66632
rect 0 65152 800 65272
rect 69200 63520 70000 63640
rect 0 62432 800 62552
rect 69200 60528 70000 60648
rect 0 59848 800 59968
rect 69200 57536 70000 57656
rect 0 57128 800 57248
rect 0 54544 800 54664
rect 69200 54680 70000 54800
rect 0 51824 800 51944
rect 69200 51688 70000 51808
rect 0 49104 800 49224
rect 69200 48696 70000 48816
rect 0 46520 800 46640
rect 69200 45704 70000 45824
rect 0 43800 800 43920
rect 69200 42712 70000 42832
rect 0 41216 800 41336
rect 69200 39856 70000 39976
rect 0 38496 800 38616
rect 69200 36864 70000 36984
rect 0 35776 800 35896
rect 69200 33872 70000 33992
rect 0 33192 800 33312
rect 69200 30880 70000 31000
rect 0 30472 800 30592
rect 0 27888 800 28008
rect 69200 28024 70000 28144
rect 0 25168 800 25288
rect 69200 25032 70000 25152
rect 0 22448 800 22568
rect 69200 22040 70000 22160
rect 0 19864 800 19984
rect 69200 19048 70000 19168
rect 0 17144 800 17264
rect 69200 16056 70000 16176
rect 0 14560 800 14680
rect 69200 13200 70000 13320
rect 0 11840 800 11960
rect 69200 10208 70000 10328
rect 0 9120 800 9240
rect 69200 7216 70000 7336
rect 0 6536 800 6656
rect 69200 4224 70000 4344
rect 0 3816 800 3936
rect 0 1232 800 1352
rect 69200 1368 70000 1488
<< obsm3 >>
rect 880 78544 69200 78573
rect 880 78400 69120 78544
rect 800 78264 69120 78400
rect 800 75960 69200 78264
rect 880 75680 69200 75960
rect 800 75552 69200 75680
rect 800 75272 69120 75552
rect 800 73376 69200 75272
rect 880 73096 69200 73376
rect 800 72560 69200 73096
rect 800 72280 69120 72560
rect 800 70656 69200 72280
rect 880 70376 69200 70656
rect 800 69568 69200 70376
rect 800 69288 69120 69568
rect 800 68072 69200 69288
rect 880 67792 69200 68072
rect 800 66712 69200 67792
rect 800 66432 69120 66712
rect 800 65352 69200 66432
rect 880 65072 69200 65352
rect 800 63720 69200 65072
rect 800 63440 69120 63720
rect 800 62632 69200 63440
rect 880 62352 69200 62632
rect 800 60728 69200 62352
rect 800 60448 69120 60728
rect 800 60048 69200 60448
rect 880 59768 69200 60048
rect 800 57736 69200 59768
rect 800 57456 69120 57736
rect 800 57328 69200 57456
rect 880 57048 69200 57328
rect 800 54880 69200 57048
rect 800 54744 69120 54880
rect 880 54600 69120 54744
rect 880 54464 69200 54600
rect 800 52024 69200 54464
rect 880 51888 69200 52024
rect 880 51744 69120 51888
rect 800 51608 69120 51744
rect 800 49304 69200 51608
rect 880 49024 69200 49304
rect 800 48896 69200 49024
rect 800 48616 69120 48896
rect 800 46720 69200 48616
rect 880 46440 69200 46720
rect 800 45904 69200 46440
rect 800 45624 69120 45904
rect 800 44000 69200 45624
rect 880 43720 69200 44000
rect 800 42912 69200 43720
rect 800 42632 69120 42912
rect 800 41416 69200 42632
rect 880 41136 69200 41416
rect 800 40056 69200 41136
rect 800 39776 69120 40056
rect 800 38696 69200 39776
rect 880 38416 69200 38696
rect 800 37064 69200 38416
rect 800 36784 69120 37064
rect 800 35976 69200 36784
rect 880 35696 69200 35976
rect 800 34072 69200 35696
rect 800 33792 69120 34072
rect 800 33392 69200 33792
rect 880 33112 69200 33392
rect 800 31080 69200 33112
rect 800 30800 69120 31080
rect 800 30672 69200 30800
rect 880 30392 69200 30672
rect 800 28224 69200 30392
rect 800 28088 69120 28224
rect 880 27944 69120 28088
rect 880 27808 69200 27944
rect 800 25368 69200 27808
rect 880 25232 69200 25368
rect 880 25088 69120 25232
rect 800 24952 69120 25088
rect 800 22648 69200 24952
rect 880 22368 69200 22648
rect 800 22240 69200 22368
rect 800 21960 69120 22240
rect 800 20064 69200 21960
rect 880 19784 69200 20064
rect 800 19248 69200 19784
rect 800 18968 69120 19248
rect 800 17344 69200 18968
rect 880 17064 69200 17344
rect 800 16256 69200 17064
rect 800 15976 69120 16256
rect 800 14760 69200 15976
rect 880 14480 69200 14760
rect 800 13400 69200 14480
rect 800 13120 69120 13400
rect 800 12040 69200 13120
rect 880 11760 69200 12040
rect 800 10408 69200 11760
rect 800 10128 69120 10408
rect 800 9320 69200 10128
rect 880 9040 69200 9320
rect 800 7416 69200 9040
rect 800 7136 69120 7416
rect 800 6736 69200 7136
rect 880 6456 69200 6736
rect 800 4424 69200 6456
rect 800 4144 69120 4424
rect 800 4016 69200 4144
rect 880 3736 69200 4016
rect 800 1568 69200 3736
rect 800 1432 69120 1568
rect 880 1288 69120 1432
rect 880 1259 69200 1288
<< metal4 >>
rect 4208 2128 4528 77840
rect 19568 2128 19888 77840
rect 34928 2128 35248 77840
rect 50288 2128 50608 77840
rect 65648 2128 65968 77840
<< obsm4 >>
rect 2083 77920 55509 78029
rect 2083 24787 4128 77920
rect 4608 24787 19488 77920
rect 19968 24787 34848 77920
rect 35328 24787 50208 77920
rect 50688 24787 55509 77920
<< labels >>
rlabel metal2 s 3882 79200 3938 80000 6 COL[0]
port 1 nsew signal input
rlabel metal2 s 6458 79200 6514 80000 6 COL[1]
port 2 nsew signal input
rlabel metal2 s 9034 79200 9090 80000 6 COL[2]
port 3 nsew signal input
rlabel metal2 s 11610 79200 11666 80000 6 COL[3]
port 4 nsew signal input
rlabel metal2 s 14186 79200 14242 80000 6 COL[4]
port 5 nsew signal input
rlabel metal3 s 69200 66512 70000 66632 6 DD[0]
port 6 nsew signal output
rlabel metal3 s 69200 69368 70000 69488 6 DD[1]
port 7 nsew signal output
rlabel metal3 s 69200 72360 70000 72480 6 DD[2]
port 8 nsew signal output
rlabel metal3 s 69200 75352 70000 75472 6 DD[3]
port 9 nsew signal output
rlabel metal3 s 69200 78344 70000 78464 6 DD[4]
port 10 nsew signal output
rlabel metal2 s 27158 79200 27214 80000 6 PWO
port 11 nsew signal input
rlabel metal2 s 29826 79200 29882 80000 6 START
port 12 nsew signal output
rlabel metal2 s 50526 79200 50582 80000 6 bcd_bus
port 13 nsew signal output
rlabel metal2 s 47950 79200 48006 80000 6 bcd_in
port 14 nsew signal input
rlabel metal2 s 53102 79200 53158 80000 6 bcd_oe
port 15 nsew signal output
rlabel metal2 s 60922 79200 60978 80000 6 carry_bus
port 16 nsew signal output
rlabel metal2 s 63498 79200 63554 80000 6 carry_in
port 17 nsew signal input
rlabel metal3 s 69200 1368 70000 1488 6 cdiv_rst
port 18 nsew signal input
rlabel metal3 s 69200 45704 70000 45824 6 dbg_arc_a1
port 19 nsew signal output
rlabel metal3 s 69200 48696 70000 48816 6 dbg_arc_b1
port 20 nsew signal output
rlabel metal3 s 69200 36864 70000 36984 6 dbg_arc_dummy
port 21 nsew signal input
rlabel metal3 s 69200 39856 70000 39976 6 dbg_arc_t1
port 22 nsew signal output
rlabel metal3 s 69200 42712 70000 42832 6 dbg_arc_t4
port 23 nsew signal output
rlabel metal3 s 69200 16056 70000 16176 6 dbg_ctc_kdn
port 24 nsew signal output
rlabel metal3 s 69200 19048 70000 19168 6 dbg_ctc_q[0]
port 25 nsew signal output
rlabel metal3 s 69200 22040 70000 22160 6 dbg_ctc_q[1]
port 26 nsew signal output
rlabel metal3 s 69200 25032 70000 25152 6 dbg_ctc_q[2]
port 27 nsew signal output
rlabel metal3 s 69200 28024 70000 28144 6 dbg_ctc_q[3]
port 28 nsew signal output
rlabel metal3 s 69200 30880 70000 31000 6 dbg_ctc_q[4]
port 29 nsew signal output
rlabel metal3 s 69200 33872 70000 33992 6 dbg_ctc_q[5]
port 30 nsew signal output
rlabel metal3 s 69200 13200 70000 13320 6 dbg_ctc_state1
port 31 nsew signal output
rlabel metal3 s 69200 51688 70000 51808 6 dbg_dsbf[0]
port 32 nsew signal output
rlabel metal3 s 69200 54680 70000 54800 6 dbg_dsbf[1]
port 33 nsew signal output
rlabel metal3 s 69200 57536 70000 57656 6 dbg_dsbf[2]
port 34 nsew signal output
rlabel metal3 s 69200 60528 70000 60648 6 dbg_dsbf[3]
port 35 nsew signal output
rlabel metal3 s 69200 63520 70000 63640 6 dbg_dsbf[4]
port 36 nsew signal output
rlabel metal2 s 62946 0 63002 800 6 dbg_enable_arc
port 37 nsew signal input
rlabel metal2 s 65798 0 65854 800 6 dbg_enable_ctc
port 38 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 dbg_enable_rom
port 39 nsew signal input
rlabel metal3 s 69200 7216 70000 7336 6 dbg_force_data
port 40 nsew signal input
rlabel metal3 s 69200 4224 70000 4344 6 dbg_internal_cdiv
port 41 nsew signal input
rlabel metal2 s 54574 0 54630 800 6 dbg_rom_roe[0]
port 42 nsew signal output
rlabel metal2 s 57334 0 57390 800 6 dbg_rom_roe[1]
port 43 nsew signal output
rlabel metal2 s 60186 0 60242 800 6 dbg_rom_roe[2]
port 44 nsew signal output
rlabel metal2 s 23754 0 23810 800 6 dbg_romdata[0]
port 45 nsew signal input
rlabel metal2 s 26514 0 26570 800 6 dbg_romdata[1]
port 46 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 dbg_romdata[2]
port 47 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 dbg_romdata[3]
port 48 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 dbg_romdata[4]
port 49 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 dbg_romdata[5]
port 50 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 dbg_romdata[6]
port 51 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 dbg_romdata[7]
port 52 nsew signal input
rlabel metal2 s 46202 0 46258 800 6 dbg_romdata[8]
port 53 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 dbg_romdata[9]
port 54 nsew signal input
rlabel metal3 s 69200 10208 70000 10328 6 dbg_sram_csb1
port 55 nsew signal input
rlabel metal2 s 58346 79200 58402 80000 6 ia_bus
port 56 nsew signal output
rlabel metal2 s 55678 79200 55734 80000 6 ia_in
port 57 nsew signal input
rlabel metal2 s 34978 79200 35034 80000 6 is_bus
port 58 nsew signal output
rlabel metal2 s 32402 79200 32458 80000 6 is_in
port 59 nsew signal input
rlabel metal2 s 37554 79200 37610 80000 6 is_oe
port 60 nsew signal output
rlabel metal2 s 1306 79200 1362 80000 6 osc_in
port 61 nsew signal input
rlabel metal2 s 16854 79200 16910 80000 6 phi1_in
port 62 nsew signal input
rlabel metal2 s 24582 79200 24638 80000 6 phi1_out
port 63 nsew signal output
rlabel metal2 s 22006 79200 22062 80000 6 phi2_in
port 64 nsew signal input
rlabel metal2 s 19430 79200 19486 80000 6 phi2_out
port 65 nsew signal output
rlabel metal2 s 1398 0 1454 800 6 sraddr_mux[0]
port 66 nsew signal output
rlabel metal2 s 4158 0 4214 800 6 sraddr_mux[1]
port 67 nsew signal output
rlabel metal2 s 6918 0 6974 800 6 sraddr_mux[2]
port 68 nsew signal output
rlabel metal2 s 9770 0 9826 800 6 sraddr_mux[3]
port 69 nsew signal output
rlabel metal2 s 12530 0 12586 800 6 sraddr_mux[4]
port 70 nsew signal output
rlabel metal2 s 15382 0 15438 800 6 sraddr_mux[5]
port 71 nsew signal output
rlabel metal2 s 18142 0 18198 800 6 sraddr_mux[6]
port 72 nsew signal output
rlabel metal2 s 20994 0 21050 800 6 sraddr_mux[7]
port 73 nsew signal output
rlabel metal2 s 51722 0 51778 800 6 sram_clk1
port 74 nsew signal output
rlabel metal3 s 0 1232 800 1352 6 srdata[0]
port 75 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 srdata[10]
port 76 nsew signal input
rlabel metal3 s 0 30472 800 30592 6 srdata[11]
port 77 nsew signal input
rlabel metal3 s 0 33192 800 33312 6 srdata[12]
port 78 nsew signal input
rlabel metal3 s 0 35776 800 35896 6 srdata[13]
port 79 nsew signal input
rlabel metal3 s 0 38496 800 38616 6 srdata[14]
port 80 nsew signal input
rlabel metal3 s 0 41216 800 41336 6 srdata[15]
port 81 nsew signal input
rlabel metal3 s 0 43800 800 43920 6 srdata[16]
port 82 nsew signal input
rlabel metal3 s 0 46520 800 46640 6 srdata[17]
port 83 nsew signal input
rlabel metal3 s 0 49104 800 49224 6 srdata[18]
port 84 nsew signal input
rlabel metal3 s 0 51824 800 51944 6 srdata[19]
port 85 nsew signal input
rlabel metal3 s 0 3816 800 3936 6 srdata[1]
port 86 nsew signal input
rlabel metal3 s 0 54544 800 54664 6 srdata[20]
port 87 nsew signal input
rlabel metal3 s 0 57128 800 57248 6 srdata[21]
port 88 nsew signal input
rlabel metal3 s 0 59848 800 59968 6 srdata[22]
port 89 nsew signal input
rlabel metal3 s 0 62432 800 62552 6 srdata[23]
port 90 nsew signal input
rlabel metal3 s 0 65152 800 65272 6 srdata[24]
port 91 nsew signal input
rlabel metal3 s 0 67872 800 67992 6 srdata[25]
port 92 nsew signal input
rlabel metal3 s 0 70456 800 70576 6 srdata[26]
port 93 nsew signal input
rlabel metal3 s 0 73176 800 73296 6 srdata[27]
port 94 nsew signal input
rlabel metal3 s 0 75760 800 75880 6 srdata[28]
port 95 nsew signal input
rlabel metal3 s 0 78480 800 78600 6 srdata[29]
port 96 nsew signal input
rlabel metal3 s 0 6536 800 6656 6 srdata[2]
port 97 nsew signal input
rlabel metal3 s 0 9120 800 9240 6 srdata[3]
port 98 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 srdata[4]
port 99 nsew signal input
rlabel metal3 s 0 14560 800 14680 6 srdata[5]
port 100 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 srdata[6]
port 101 nsew signal input
rlabel metal3 s 0 19864 800 19984 6 srdata[7]
port 102 nsew signal input
rlabel metal3 s 0 22448 800 22568 6 srdata[8]
port 103 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 srdata[9]
port 104 nsew signal input
rlabel metal2 s 66074 79200 66130 80000 6 sync_bus
port 105 nsew signal output
rlabel metal2 s 68650 79200 68706 80000 6 sync_in
port 106 nsew signal input
rlabel metal4 s 4208 2128 4528 77840 6 vccd1
port 107 nsew power input
rlabel metal4 s 34928 2128 35248 77840 6 vccd1
port 107 nsew power input
rlabel metal4 s 65648 2128 65968 77840 6 vccd1
port 107 nsew power input
rlabel metal4 s 19568 2128 19888 77840 6 vssd1
port 108 nsew ground input
rlabel metal4 s 50288 2128 50608 77840 6 vssd1
port 108 nsew ground input
rlabel metal2 s 42706 79200 42762 80000 6 ws_bus
port 109 nsew signal output
rlabel metal2 s 40130 79200 40186 80000 6 ws_in
port 110 nsew signal input
rlabel metal2 s 45374 79200 45430 80000 6 ws_oe
port 111 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 70000 80000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9124676
string GDS_FILE /home/andylithia/openmpw/MPWTRIAL/openlane/hp35_core/runs/hp35_core/results/finishing/hp35_core.magic.gds
string GDS_START 1145738
<< end >>

