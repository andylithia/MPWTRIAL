VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO hp35_core
  CLASS BLOCK ;
  FOREIGN hp35_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 350.000 BY 400.000 ;
  PIN COL[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 396.000 16.930 400.000 ;
    END
  END COL[0]
  PIN COL[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 396.000 28.430 400.000 ;
    END
  END COL[1]
  PIN COL[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 396.000 39.470 400.000 ;
    END
  END COL[2]
  PIN COL[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 396.000 50.970 400.000 ;
    END
  END COL[3]
  PIN COL[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 396.000 62.010 400.000 ;
    END
  END COL[4]
  PIN DD[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 332.560 350.000 333.160 ;
    END
  END DD[0]
  PIN DD[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 346.840 350.000 347.440 ;
    END
  END DD[1]
  PIN DD[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 361.800 350.000 362.400 ;
    END
  END DD[2]
  PIN DD[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 376.760 350.000 377.360 ;
    END
  END DD[3]
  PIN DD[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 391.720 350.000 392.320 ;
    END
  END DD[4]
  PIN PWO
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 396.000 130.090 400.000 ;
    END
  END PWO
  PIN START
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 396.000 141.130 400.000 ;
    END
  END START
  PIN bcd_bus
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 396.000 231.290 400.000 ;
    END
  END bcd_bus
  PIN bcd_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 396.000 220.250 400.000 ;
    END
  END bcd_in
  PIN bcd_oen
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 396.000 242.790 400.000 ;
    END
  END bcd_oen
  PIN carry_bus
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 396.000 287.870 400.000 ;
    END
  END carry_bus
  PIN carry_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.090 396.000 299.370 400.000 ;
    END
  END carry_in
  PIN carry_oen
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.130 396.000 310.410 400.000 ;
    END
  END carry_oen
  PIN cdiv_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 6.840 350.000 7.440 ;
    END
  END cdiv_rst
  PIN dbg_arc_a1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 228.520 350.000 229.120 ;
    END
  END dbg_arc_a1
  PIN dbg_arc_b1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 243.480 350.000 244.080 ;
    END
  END dbg_arc_b1
  PIN dbg_arc_dummy
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 184.320 350.000 184.920 ;
    END
  END dbg_arc_dummy
  PIN dbg_arc_t1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 199.280 350.000 199.880 ;
    END
  END dbg_arc_t1
  PIN dbg_arc_t4
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 213.560 350.000 214.160 ;
    END
  END dbg_arc_t4
  PIN dbg_ctc_kdn
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 80.280 350.000 80.880 ;
    END
  END dbg_ctc_kdn
  PIN dbg_ctc_q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 95.240 350.000 95.840 ;
    END
  END dbg_ctc_q[0]
  PIN dbg_ctc_q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 110.200 350.000 110.800 ;
    END
  END dbg_ctc_q[1]
  PIN dbg_ctc_q[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 125.160 350.000 125.760 ;
    END
  END dbg_ctc_q[2]
  PIN dbg_ctc_q[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 140.120 350.000 140.720 ;
    END
  END dbg_ctc_q[3]
  PIN dbg_ctc_q[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 154.400 350.000 155.000 ;
    END
  END dbg_ctc_q[4]
  PIN dbg_ctc_q[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 169.360 350.000 169.960 ;
    END
  END dbg_ctc_q[5]
  PIN dbg_ctc_state1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 66.000 350.000 66.600 ;
    END
  END dbg_ctc_state1
  PIN dbg_disable_arc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 0.000 315.010 4.000 ;
    END
  END dbg_disable_arc
  PIN dbg_disable_ctc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.990 0.000 329.270 4.000 ;
    END
  END dbg_disable_ctc
  PIN dbg_disable_rom
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 0.000 343.070 4.000 ;
    END
  END dbg_disable_rom
  PIN dbg_dsbf[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 258.440 350.000 259.040 ;
    END
  END dbg_dsbf[0]
  PIN dbg_dsbf[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 273.400 350.000 274.000 ;
    END
  END dbg_dsbf[1]
  PIN dbg_dsbf[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 287.680 350.000 288.280 ;
    END
  END dbg_dsbf[2]
  PIN dbg_dsbf[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 302.640 350.000 303.240 ;
    END
  END dbg_dsbf[3]
  PIN dbg_dsbf[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 317.600 350.000 318.200 ;
    END
  END dbg_dsbf[4]
  PIN dbg_force_data
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 36.080 350.000 36.680 ;
    END
  END dbg_force_data
  PIN dbg_internal_cdiv
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 21.120 350.000 21.720 ;
    END
  END dbg_internal_cdiv
  PIN dbg_rom_roe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 0.000 273.150 4.000 ;
    END
  END dbg_rom_roe[0]
  PIN dbg_rom_roe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END dbg_rom_roe[1]
  PIN dbg_rom_roe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 0.000 301.210 4.000 ;
    END
  END dbg_rom_roe[2]
  PIN dbg_romdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END dbg_romdata[0]
  PIN dbg_romdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 4.000 ;
    END
  END dbg_romdata[1]
  PIN dbg_romdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 4.000 ;
    END
  END dbg_romdata[2]
  PIN dbg_romdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 4.000 ;
    END
  END dbg_romdata[3]
  PIN dbg_romdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END dbg_romdata[4]
  PIN dbg_romdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 0.000 188.970 4.000 ;
    END
  END dbg_romdata[5]
  PIN dbg_romdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END dbg_romdata[6]
  PIN dbg_romdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 0.000 217.030 4.000 ;
    END
  END dbg_romdata[7]
  PIN dbg_romdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END dbg_romdata[8]
  PIN dbg_romdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END dbg_romdata[9]
  PIN dbg_sram_csb1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 51.040 350.000 51.640 ;
    END
  END dbg_sram_csb1
  PIN ia_bus
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 396.000 265.330 400.000 ;
    END
  END ia_bus
  PIN ia_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 396.000 254.290 400.000 ;
    END
  END ia_in
  PIN ia_oen
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.550 396.000 276.830 400.000 ;
    END
  END ia_oen
  PIN is_bus
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 396.000 163.670 400.000 ;
    END
  END is_bus
  PIN is_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 396.000 152.630 400.000 ;
    END
  END is_in
  PIN is_oen
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 396.000 175.170 400.000 ;
    END
  END is_oen
  PIN osc_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 396.000 5.890 400.000 ;
    END
  END osc_in
  PIN phi1_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 396.000 73.510 400.000 ;
    END
  END phi1_in
  PIN phi1_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 396.000 107.090 400.000 ;
    END
  END phi1_out
  PIN phi2_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 396.000 96.050 400.000 ;
    END
  END phi2_in
  PIN phi2_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 396.000 84.550 400.000 ;
    END
  END phi2_out
  PIN phi_oen
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 396.000 118.590 400.000 ;
    END
  END phi_oen
  PIN sraddr_mux[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END sraddr_mux[0]
  PIN sraddr_mux[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END sraddr_mux[1]
  PIN sraddr_mux[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 4.000 ;
    END
  END sraddr_mux[2]
  PIN sraddr_mux[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END sraddr_mux[3]
  PIN sraddr_mux[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END sraddr_mux[4]
  PIN sraddr_mux[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 4.000 ;
    END
  END sraddr_mux[5]
  PIN sraddr_mux[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 0.000 90.990 4.000 ;
    END
  END sraddr_mux[6]
  PIN sraddr_mux[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 4.000 ;
    END
  END sraddr_mux[7]
  PIN sram_clk1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END sram_clk1
  PIN srdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.160 4.000 6.760 ;
    END
  END srdata[0]
  PIN srdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END srdata[10]
  PIN srdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END srdata[11]
  PIN srdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END srdata[12]
  PIN srdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.880 4.000 179.480 ;
    END
  END srdata[13]
  PIN srdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 192.480 4.000 193.080 ;
    END
  END srdata[14]
  PIN srdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.080 4.000 206.680 ;
    END
  END srdata[15]
  PIN srdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.000 4.000 219.600 ;
    END
  END srdata[16]
  PIN srdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END srdata[17]
  PIN srdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 245.520 4.000 246.120 ;
    END
  END srdata[18]
  PIN srdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.120 4.000 259.720 ;
    END
  END srdata[19]
  PIN srdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END srdata[1]
  PIN srdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.720 4.000 273.320 ;
    END
  END srdata[20]
  PIN srdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END srdata[21]
  PIN srdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END srdata[22]
  PIN srdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.160 4.000 312.760 ;
    END
  END srdata[23]
  PIN srdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.760 4.000 326.360 ;
    END
  END srdata[24]
  PIN srdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 339.360 4.000 339.960 ;
    END
  END srdata[25]
  PIN srdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.280 4.000 352.880 ;
    END
  END srdata[26]
  PIN srdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.880 4.000 366.480 ;
    END
  END srdata[27]
  PIN srdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.800 4.000 379.400 ;
    END
  END srdata[28]
  PIN srdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 392.400 4.000 393.000 ;
    END
  END srdata[29]
  PIN srdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END srdata[2]
  PIN srdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 4.000 46.200 ;
    END
  END srdata[3]
  PIN srdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 4.000 59.800 ;
    END
  END srdata[4]
  PIN srdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 4.000 73.400 ;
    END
  END srdata[5]
  PIN srdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END srdata[6]
  PIN srdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END srdata[7]
  PIN srdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END srdata[8]
  PIN srdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END srdata[9]
  PIN sync_bus
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 396.000 321.910 400.000 ;
    END
  END sync_bus
  PIN sync_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 396.000 332.950 400.000 ;
    END
  END sync_in
  PIN sync_oen
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 396.000 344.450 400.000 ;
    END
  END sync_oen
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 389.200 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 389.200 ;
    END
  END vssd1
  PIN ws_bus
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 396.000 197.710 400.000 ;
    END
  END ws_bus
  PIN ws_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 396.000 186.210 400.000 ;
    END
  END ws_in
  PIN ws_oen
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 396.000 208.750 400.000 ;
    END
  END ws_oen
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 344.080 389.045 ;
      LAYER met1 ;
        RECT 5.520 9.220 344.470 389.200 ;
      LAYER met2 ;
        RECT 6.170 395.720 16.370 396.000 ;
        RECT 17.210 395.720 27.870 396.000 ;
        RECT 28.710 395.720 38.910 396.000 ;
        RECT 39.750 395.720 50.410 396.000 ;
        RECT 51.250 395.720 61.450 396.000 ;
        RECT 62.290 395.720 72.950 396.000 ;
        RECT 73.790 395.720 83.990 396.000 ;
        RECT 84.830 395.720 95.490 396.000 ;
        RECT 96.330 395.720 106.530 396.000 ;
        RECT 107.370 395.720 118.030 396.000 ;
        RECT 118.870 395.720 129.530 396.000 ;
        RECT 130.370 395.720 140.570 396.000 ;
        RECT 141.410 395.720 152.070 396.000 ;
        RECT 152.910 395.720 163.110 396.000 ;
        RECT 163.950 395.720 174.610 396.000 ;
        RECT 175.450 395.720 185.650 396.000 ;
        RECT 186.490 395.720 197.150 396.000 ;
        RECT 197.990 395.720 208.190 396.000 ;
        RECT 209.030 395.720 219.690 396.000 ;
        RECT 220.530 395.720 230.730 396.000 ;
        RECT 231.570 395.720 242.230 396.000 ;
        RECT 243.070 395.720 253.730 396.000 ;
        RECT 254.570 395.720 264.770 396.000 ;
        RECT 265.610 395.720 276.270 396.000 ;
        RECT 277.110 395.720 287.310 396.000 ;
        RECT 288.150 395.720 298.810 396.000 ;
        RECT 299.650 395.720 309.850 396.000 ;
        RECT 310.690 395.720 321.350 396.000 ;
        RECT 322.190 395.720 332.390 396.000 ;
        RECT 333.230 395.720 343.890 396.000 ;
        RECT 5.620 4.280 344.440 395.720 ;
        RECT 5.620 4.000 6.710 4.280 ;
        RECT 7.550 4.000 20.510 4.280 ;
        RECT 21.350 4.000 34.310 4.280 ;
        RECT 35.150 4.000 48.570 4.280 ;
        RECT 49.410 4.000 62.370 4.280 ;
        RECT 63.210 4.000 76.630 4.280 ;
        RECT 77.470 4.000 90.430 4.280 ;
        RECT 91.270 4.000 104.690 4.280 ;
        RECT 105.530 4.000 118.490 4.280 ;
        RECT 119.330 4.000 132.290 4.280 ;
        RECT 133.130 4.000 146.550 4.280 ;
        RECT 147.390 4.000 160.350 4.280 ;
        RECT 161.190 4.000 174.610 4.280 ;
        RECT 175.450 4.000 188.410 4.280 ;
        RECT 189.250 4.000 202.670 4.280 ;
        RECT 203.510 4.000 216.470 4.280 ;
        RECT 217.310 4.000 230.730 4.280 ;
        RECT 231.570 4.000 244.530 4.280 ;
        RECT 245.370 4.000 258.330 4.280 ;
        RECT 259.170 4.000 272.590 4.280 ;
        RECT 273.430 4.000 286.390 4.280 ;
        RECT 287.230 4.000 300.650 4.280 ;
        RECT 301.490 4.000 314.450 4.280 ;
        RECT 315.290 4.000 328.710 4.280 ;
        RECT 329.550 4.000 342.510 4.280 ;
        RECT 343.350 4.000 344.440 4.280 ;
      LAYER met3 ;
        RECT 4.400 392.720 346.000 392.865 ;
        RECT 4.400 392.000 345.600 392.720 ;
        RECT 4.000 391.320 345.600 392.000 ;
        RECT 4.000 379.800 346.000 391.320 ;
        RECT 4.400 378.400 346.000 379.800 ;
        RECT 4.000 377.760 346.000 378.400 ;
        RECT 4.000 376.360 345.600 377.760 ;
        RECT 4.000 366.880 346.000 376.360 ;
        RECT 4.400 365.480 346.000 366.880 ;
        RECT 4.000 362.800 346.000 365.480 ;
        RECT 4.000 361.400 345.600 362.800 ;
        RECT 4.000 353.280 346.000 361.400 ;
        RECT 4.400 351.880 346.000 353.280 ;
        RECT 4.000 347.840 346.000 351.880 ;
        RECT 4.000 346.440 345.600 347.840 ;
        RECT 4.000 340.360 346.000 346.440 ;
        RECT 4.400 338.960 346.000 340.360 ;
        RECT 4.000 333.560 346.000 338.960 ;
        RECT 4.000 332.160 345.600 333.560 ;
        RECT 4.000 326.760 346.000 332.160 ;
        RECT 4.400 325.360 346.000 326.760 ;
        RECT 4.000 318.600 346.000 325.360 ;
        RECT 4.000 317.200 345.600 318.600 ;
        RECT 4.000 313.160 346.000 317.200 ;
        RECT 4.400 311.760 346.000 313.160 ;
        RECT 4.000 303.640 346.000 311.760 ;
        RECT 4.000 302.240 345.600 303.640 ;
        RECT 4.000 300.240 346.000 302.240 ;
        RECT 4.400 298.840 346.000 300.240 ;
        RECT 4.000 288.680 346.000 298.840 ;
        RECT 4.000 287.280 345.600 288.680 ;
        RECT 4.000 286.640 346.000 287.280 ;
        RECT 4.400 285.240 346.000 286.640 ;
        RECT 4.000 274.400 346.000 285.240 ;
        RECT 4.000 273.720 345.600 274.400 ;
        RECT 4.400 273.000 345.600 273.720 ;
        RECT 4.400 272.320 346.000 273.000 ;
        RECT 4.000 260.120 346.000 272.320 ;
        RECT 4.400 259.440 346.000 260.120 ;
        RECT 4.400 258.720 345.600 259.440 ;
        RECT 4.000 258.040 345.600 258.720 ;
        RECT 4.000 246.520 346.000 258.040 ;
        RECT 4.400 245.120 346.000 246.520 ;
        RECT 4.000 244.480 346.000 245.120 ;
        RECT 4.000 243.080 345.600 244.480 ;
        RECT 4.000 233.600 346.000 243.080 ;
        RECT 4.400 232.200 346.000 233.600 ;
        RECT 4.000 229.520 346.000 232.200 ;
        RECT 4.000 228.120 345.600 229.520 ;
        RECT 4.000 220.000 346.000 228.120 ;
        RECT 4.400 218.600 346.000 220.000 ;
        RECT 4.000 214.560 346.000 218.600 ;
        RECT 4.000 213.160 345.600 214.560 ;
        RECT 4.000 207.080 346.000 213.160 ;
        RECT 4.400 205.680 346.000 207.080 ;
        RECT 4.000 200.280 346.000 205.680 ;
        RECT 4.000 198.880 345.600 200.280 ;
        RECT 4.000 193.480 346.000 198.880 ;
        RECT 4.400 192.080 346.000 193.480 ;
        RECT 4.000 185.320 346.000 192.080 ;
        RECT 4.000 183.920 345.600 185.320 ;
        RECT 4.000 179.880 346.000 183.920 ;
        RECT 4.400 178.480 346.000 179.880 ;
        RECT 4.000 170.360 346.000 178.480 ;
        RECT 4.000 168.960 345.600 170.360 ;
        RECT 4.000 166.960 346.000 168.960 ;
        RECT 4.400 165.560 346.000 166.960 ;
        RECT 4.000 155.400 346.000 165.560 ;
        RECT 4.000 154.000 345.600 155.400 ;
        RECT 4.000 153.360 346.000 154.000 ;
        RECT 4.400 151.960 346.000 153.360 ;
        RECT 4.000 141.120 346.000 151.960 ;
        RECT 4.000 140.440 345.600 141.120 ;
        RECT 4.400 139.720 345.600 140.440 ;
        RECT 4.400 139.040 346.000 139.720 ;
        RECT 4.000 126.840 346.000 139.040 ;
        RECT 4.400 126.160 346.000 126.840 ;
        RECT 4.400 125.440 345.600 126.160 ;
        RECT 4.000 124.760 345.600 125.440 ;
        RECT 4.000 113.240 346.000 124.760 ;
        RECT 4.400 111.840 346.000 113.240 ;
        RECT 4.000 111.200 346.000 111.840 ;
        RECT 4.000 109.800 345.600 111.200 ;
        RECT 4.000 100.320 346.000 109.800 ;
        RECT 4.400 98.920 346.000 100.320 ;
        RECT 4.000 96.240 346.000 98.920 ;
        RECT 4.000 94.840 345.600 96.240 ;
        RECT 4.000 86.720 346.000 94.840 ;
        RECT 4.400 85.320 346.000 86.720 ;
        RECT 4.000 81.280 346.000 85.320 ;
        RECT 4.000 79.880 345.600 81.280 ;
        RECT 4.000 73.800 346.000 79.880 ;
        RECT 4.400 72.400 346.000 73.800 ;
        RECT 4.000 67.000 346.000 72.400 ;
        RECT 4.000 65.600 345.600 67.000 ;
        RECT 4.000 60.200 346.000 65.600 ;
        RECT 4.400 58.800 346.000 60.200 ;
        RECT 4.000 52.040 346.000 58.800 ;
        RECT 4.000 50.640 345.600 52.040 ;
        RECT 4.000 46.600 346.000 50.640 ;
        RECT 4.400 45.200 346.000 46.600 ;
        RECT 4.000 37.080 346.000 45.200 ;
        RECT 4.000 35.680 345.600 37.080 ;
        RECT 4.000 33.680 346.000 35.680 ;
        RECT 4.400 32.280 346.000 33.680 ;
        RECT 4.000 22.120 346.000 32.280 ;
        RECT 4.000 20.720 345.600 22.120 ;
        RECT 4.000 20.080 346.000 20.720 ;
        RECT 4.400 18.680 346.000 20.080 ;
        RECT 4.000 7.840 346.000 18.680 ;
        RECT 4.000 7.160 345.600 7.840 ;
        RECT 4.400 6.440 345.600 7.160 ;
        RECT 4.400 6.295 346.000 6.440 ;
      LAYER met4 ;
        RECT 8.575 93.335 20.640 386.745 ;
        RECT 23.040 93.335 97.440 386.745 ;
        RECT 99.840 93.335 174.240 386.745 ;
        RECT 176.640 93.335 251.040 386.745 ;
        RECT 253.440 93.335 268.345 386.745 ;
  END
END hp35_core
END LIBRARY

