magic
tech sky130A
magscale 1 2
timestamp 1654387249
<< obsli1 >>
rect 1104 2159 98808 297585
<< obsm1 >>
rect 1104 2128 98808 297616
<< metal2 >>
rect 1490 299200 1546 300000
rect 4526 299200 4582 300000
rect 7654 299200 7710 300000
rect 10782 299200 10838 300000
rect 13910 299200 13966 300000
rect 17038 299200 17094 300000
rect 20166 299200 20222 300000
rect 23294 299200 23350 300000
rect 26422 299200 26478 300000
rect 29550 299200 29606 300000
rect 32678 299200 32734 300000
rect 35806 299200 35862 300000
rect 38934 299200 38990 300000
rect 42062 299200 42118 300000
rect 45190 299200 45246 300000
rect 48318 299200 48374 300000
rect 51446 299200 51502 300000
rect 54574 299200 54630 300000
rect 57702 299200 57758 300000
rect 60830 299200 60886 300000
rect 63958 299200 64014 300000
rect 67086 299200 67142 300000
rect 70214 299200 70270 300000
rect 73342 299200 73398 300000
rect 76470 299200 76526 300000
rect 79598 299200 79654 300000
rect 82726 299200 82782 300000
rect 85854 299200 85910 300000
rect 88982 299200 89038 300000
rect 92110 299200 92166 300000
rect 95238 299200 95294 300000
rect 98366 299200 98422 300000
rect 2778 0 2834 800
rect 8298 0 8354 800
rect 13818 0 13874 800
rect 19430 0 19486 800
rect 24950 0 25006 800
rect 30470 0 30526 800
rect 36082 0 36138 800
rect 41602 0 41658 800
rect 47214 0 47270 800
rect 52734 0 52790 800
rect 58254 0 58310 800
rect 63866 0 63922 800
rect 69386 0 69442 800
rect 74998 0 75054 800
rect 80518 0 80574 800
rect 86038 0 86094 800
rect 91650 0 91706 800
rect 97170 0 97226 800
<< obsm2 >>
rect 1398 299144 1434 299200
rect 1602 299144 4470 299200
rect 4638 299144 7598 299200
rect 7766 299144 10726 299200
rect 10894 299144 13854 299200
rect 14022 299144 16982 299200
rect 17150 299144 20110 299200
rect 20278 299144 23238 299200
rect 23406 299144 26366 299200
rect 26534 299144 29494 299200
rect 29662 299144 32622 299200
rect 32790 299144 35750 299200
rect 35918 299144 38878 299200
rect 39046 299144 42006 299200
rect 42174 299144 45134 299200
rect 45302 299144 48262 299200
rect 48430 299144 51390 299200
rect 51558 299144 54518 299200
rect 54686 299144 57646 299200
rect 57814 299144 60774 299200
rect 60942 299144 63902 299200
rect 64070 299144 67030 299200
rect 67198 299144 70158 299200
rect 70326 299144 73286 299200
rect 73454 299144 76414 299200
rect 76582 299144 79542 299200
rect 79710 299144 82670 299200
rect 82838 299144 85798 299200
rect 85966 299144 88926 299200
rect 89094 299144 92054 299200
rect 92222 299144 95182 299200
rect 95350 299144 98310 299200
rect 98478 299144 98514 299200
rect 1398 856 98514 299144
rect 1398 800 2722 856
rect 2890 800 8242 856
rect 8410 800 13762 856
rect 13930 800 19374 856
rect 19542 800 24894 856
rect 25062 800 30414 856
rect 30582 800 36026 856
rect 36194 800 41546 856
rect 41714 800 47158 856
rect 47326 800 52678 856
rect 52846 800 58198 856
rect 58366 800 63810 856
rect 63978 800 69330 856
rect 69498 800 74942 856
rect 75110 800 80462 856
rect 80630 800 85982 856
rect 86150 800 91594 856
rect 91762 800 97114 856
rect 97282 800 98514 856
<< metal3 >>
rect 0 296216 800 296336
rect 99200 292408 100000 292528
rect 0 288872 800 288992
rect 0 281528 800 281648
rect 99200 277448 100000 277568
rect 0 274184 800 274304
rect 0 266840 800 266960
rect 99200 262488 100000 262608
rect 0 259632 800 259752
rect 0 252288 800 252408
rect 99200 247392 100000 247512
rect 0 244944 800 245064
rect 0 237600 800 237720
rect 99200 232432 100000 232552
rect 0 230256 800 230376
rect 0 223048 800 223168
rect 99200 217472 100000 217592
rect 0 215704 800 215824
rect 0 208360 800 208480
rect 99200 202376 100000 202496
rect 0 201016 800 201136
rect 0 193672 800 193792
rect 99200 187416 100000 187536
rect 0 186464 800 186584
rect 0 179120 800 179240
rect 99200 172456 100000 172576
rect 0 171776 800 171896
rect 0 164432 800 164552
rect 99200 157496 100000 157616
rect 0 157088 800 157208
rect 0 149880 800 150000
rect 0 142536 800 142656
rect 99200 142400 100000 142520
rect 0 135192 800 135312
rect 0 127848 800 127968
rect 99200 127440 100000 127560
rect 0 120504 800 120624
rect 0 113296 800 113416
rect 99200 112480 100000 112600
rect 0 105952 800 106072
rect 0 98608 800 98728
rect 99200 97384 100000 97504
rect 0 91264 800 91384
rect 0 83920 800 84040
rect 99200 82424 100000 82544
rect 0 76712 800 76832
rect 0 69368 800 69488
rect 99200 67464 100000 67584
rect 0 62024 800 62144
rect 0 54680 800 54800
rect 99200 52368 100000 52488
rect 0 47336 800 47456
rect 0 40128 800 40248
rect 99200 37408 100000 37528
rect 0 32784 800 32904
rect 0 25440 800 25560
rect 99200 22448 100000 22568
rect 0 18096 800 18216
rect 0 10752 800 10872
rect 99200 7488 100000 7608
rect 0 3544 800 3664
<< obsm3 >>
rect 800 296416 99200 297601
rect 880 296136 99200 296416
rect 800 292608 99200 296136
rect 800 292328 99120 292608
rect 800 289072 99200 292328
rect 880 288792 99200 289072
rect 800 281728 99200 288792
rect 880 281448 99200 281728
rect 800 277648 99200 281448
rect 800 277368 99120 277648
rect 800 274384 99200 277368
rect 880 274104 99200 274384
rect 800 267040 99200 274104
rect 880 266760 99200 267040
rect 800 262688 99200 266760
rect 800 262408 99120 262688
rect 800 259832 99200 262408
rect 880 259552 99200 259832
rect 800 252488 99200 259552
rect 880 252208 99200 252488
rect 800 247592 99200 252208
rect 800 247312 99120 247592
rect 800 245144 99200 247312
rect 880 244864 99200 245144
rect 800 237800 99200 244864
rect 880 237520 99200 237800
rect 800 232632 99200 237520
rect 800 232352 99120 232632
rect 800 230456 99200 232352
rect 880 230176 99200 230456
rect 800 223248 99200 230176
rect 880 222968 99200 223248
rect 800 217672 99200 222968
rect 800 217392 99120 217672
rect 800 215904 99200 217392
rect 880 215624 99200 215904
rect 800 208560 99200 215624
rect 880 208280 99200 208560
rect 800 202576 99200 208280
rect 800 202296 99120 202576
rect 800 201216 99200 202296
rect 880 200936 99200 201216
rect 800 193872 99200 200936
rect 880 193592 99200 193872
rect 800 187616 99200 193592
rect 800 187336 99120 187616
rect 800 186664 99200 187336
rect 880 186384 99200 186664
rect 800 179320 99200 186384
rect 880 179040 99200 179320
rect 800 172656 99200 179040
rect 800 172376 99120 172656
rect 800 171976 99200 172376
rect 880 171696 99200 171976
rect 800 164632 99200 171696
rect 880 164352 99200 164632
rect 800 157696 99200 164352
rect 800 157416 99120 157696
rect 800 157288 99200 157416
rect 880 157008 99200 157288
rect 800 150080 99200 157008
rect 880 149800 99200 150080
rect 800 142736 99200 149800
rect 880 142600 99200 142736
rect 880 142456 99120 142600
rect 800 142320 99120 142456
rect 800 135392 99200 142320
rect 880 135112 99200 135392
rect 800 128048 99200 135112
rect 880 127768 99200 128048
rect 800 127640 99200 127768
rect 800 127360 99120 127640
rect 800 120704 99200 127360
rect 880 120424 99200 120704
rect 800 113496 99200 120424
rect 880 113216 99200 113496
rect 800 112680 99200 113216
rect 800 112400 99120 112680
rect 800 106152 99200 112400
rect 880 105872 99200 106152
rect 800 98808 99200 105872
rect 880 98528 99200 98808
rect 800 97584 99200 98528
rect 800 97304 99120 97584
rect 800 91464 99200 97304
rect 880 91184 99200 91464
rect 800 84120 99200 91184
rect 880 83840 99200 84120
rect 800 82624 99200 83840
rect 800 82344 99120 82624
rect 800 76912 99200 82344
rect 880 76632 99200 76912
rect 800 69568 99200 76632
rect 880 69288 99200 69568
rect 800 67664 99200 69288
rect 800 67384 99120 67664
rect 800 62224 99200 67384
rect 880 61944 99200 62224
rect 800 54880 99200 61944
rect 880 54600 99200 54880
rect 800 52568 99200 54600
rect 800 52288 99120 52568
rect 800 47536 99200 52288
rect 880 47256 99200 47536
rect 800 40328 99200 47256
rect 880 40048 99200 40328
rect 800 37608 99200 40048
rect 800 37328 99120 37608
rect 800 32984 99200 37328
rect 880 32704 99200 32984
rect 800 25640 99200 32704
rect 880 25360 99200 25640
rect 800 22648 99200 25360
rect 800 22368 99120 22648
rect 800 18296 99200 22368
rect 880 18016 99200 18296
rect 800 10952 99200 18016
rect 880 10672 99200 10952
rect 800 7688 99200 10672
rect 800 7408 99120 7688
rect 800 3744 99200 7408
rect 880 3464 99200 3744
rect 800 2143 99200 3464
<< metal4 >>
rect 4208 2128 4528 297616
rect 19568 2128 19888 297616
rect 34928 2128 35248 297616
rect 50288 2128 50608 297616
rect 65648 2128 65968 297616
rect 81008 2128 81328 297616
rect 96368 2128 96688 297616
<< obsm4 >>
rect 24531 2619 34848 297125
rect 35328 2619 50208 297125
rect 50688 2619 64893 297125
<< labels >>
rlabel metal2 s 4526 299200 4582 300000 6 COL[0]
port 1 nsew signal input
rlabel metal2 s 7654 299200 7710 300000 6 COL[1]
port 2 nsew signal input
rlabel metal2 s 10782 299200 10838 300000 6 COL[2]
port 3 nsew signal input
rlabel metal2 s 13910 299200 13966 300000 6 COL[3]
port 4 nsew signal input
rlabel metal2 s 17038 299200 17094 300000 6 COL[4]
port 5 nsew signal input
rlabel metal2 s 35806 299200 35862 300000 6 DD[0]
port 6 nsew signal output
rlabel metal2 s 38934 299200 38990 300000 6 DD[1]
port 7 nsew signal output
rlabel metal2 s 42062 299200 42118 300000 6 DD[2]
port 8 nsew signal output
rlabel metal2 s 45190 299200 45246 300000 6 DD[3]
port 9 nsew signal output
rlabel metal2 s 48318 299200 48374 300000 6 DD[4]
port 10 nsew signal output
rlabel metal2 s 32678 299200 32734 300000 6 PWO
port 11 nsew signal input
rlabel metal2 s 51446 299200 51502 300000 6 START
port 12 nsew signal output
rlabel metal2 s 76470 299200 76526 300000 6 bcd_bus
port 13 nsew signal output
rlabel metal2 s 73342 299200 73398 300000 6 bcd_in
port 14 nsew signal input
rlabel metal2 s 79598 299200 79654 300000 6 bcd_oe
port 15 nsew signal output
rlabel metal2 s 88982 299200 89038 300000 6 carry_bus
port 16 nsew signal output
rlabel metal2 s 92110 299200 92166 300000 6 carry_in
port 17 nsew signal input
rlabel metal3 s 99200 7488 100000 7608 6 cdiv_rst
port 18 nsew signal input
rlabel metal2 s 47214 0 47270 800 6 dbg_arc_a1
port 19 nsew signal output
rlabel metal2 s 52734 0 52790 800 6 dbg_arc_b1
port 20 nsew signal output
rlabel metal2 s 19430 0 19486 800 6 dbg_arc_dummy
port 21 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 dbg_arc_t1
port 22 nsew signal output
rlabel metal2 s 41602 0 41658 800 6 dbg_arc_t4
port 23 nsew signal output
rlabel metal2 s 63866 0 63922 800 6 dbg_ctc_kdn
port 24 nsew signal output
rlabel metal2 s 69386 0 69442 800 6 dbg_ctc_q[0]
port 25 nsew signal output
rlabel metal2 s 74998 0 75054 800 6 dbg_ctc_q[1]
port 26 nsew signal output
rlabel metal2 s 80518 0 80574 800 6 dbg_ctc_q[2]
port 27 nsew signal output
rlabel metal2 s 86038 0 86094 800 6 dbg_ctc_q[3]
port 28 nsew signal output
rlabel metal2 s 91650 0 91706 800 6 dbg_ctc_q[4]
port 29 nsew signal output
rlabel metal2 s 97170 0 97226 800 6 dbg_ctc_q[5]
port 30 nsew signal output
rlabel metal2 s 58254 0 58310 800 6 dbg_ctc_state1
port 31 nsew signal output
rlabel metal3 s 99200 232432 100000 232552 6 dbg_dsbf[0]
port 32 nsew signal output
rlabel metal3 s 99200 247392 100000 247512 6 dbg_dsbf[1]
port 33 nsew signal output
rlabel metal3 s 99200 262488 100000 262608 6 dbg_dsbf[2]
port 34 nsew signal output
rlabel metal3 s 99200 277448 100000 277568 6 dbg_dsbf[3]
port 35 nsew signal output
rlabel metal3 s 99200 292408 100000 292528 6 dbg_dsbf[4]
port 36 nsew signal output
rlabel metal2 s 2778 0 2834 800 6 dbg_enable_arc
port 37 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 dbg_enable_ctc
port 38 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 dbg_enable_rom
port 39 nsew signal input
rlabel metal2 s 24950 0 25006 800 6 dbg_force_data
port 40 nsew signal input
rlabel metal3 s 99200 22448 100000 22568 6 dbg_internal_cdiv
port 41 nsew signal input
rlabel metal3 s 99200 187416 100000 187536 6 dbg_rom_roe[0]
port 42 nsew signal output
rlabel metal3 s 99200 202376 100000 202496 6 dbg_rom_roe[1]
port 43 nsew signal output
rlabel metal3 s 99200 217472 100000 217592 6 dbg_rom_roe[2]
port 44 nsew signal output
rlabel metal3 s 99200 37408 100000 37528 6 dbg_romdata[0]
port 45 nsew signal input
rlabel metal3 s 99200 52368 100000 52488 6 dbg_romdata[1]
port 46 nsew signal input
rlabel metal3 s 99200 67464 100000 67584 6 dbg_romdata[2]
port 47 nsew signal input
rlabel metal3 s 99200 82424 100000 82544 6 dbg_romdata[3]
port 48 nsew signal input
rlabel metal3 s 99200 97384 100000 97504 6 dbg_romdata[4]
port 49 nsew signal input
rlabel metal3 s 99200 112480 100000 112600 6 dbg_romdata[5]
port 50 nsew signal input
rlabel metal3 s 99200 127440 100000 127560 6 dbg_romdata[6]
port 51 nsew signal input
rlabel metal3 s 99200 142400 100000 142520 6 dbg_romdata[7]
port 52 nsew signal input
rlabel metal3 s 99200 157496 100000 157616 6 dbg_romdata[8]
port 53 nsew signal input
rlabel metal3 s 99200 172456 100000 172576 6 dbg_romdata[9]
port 54 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 dbg_sram_csb1
port 55 nsew signal input
rlabel metal2 s 85854 299200 85910 300000 6 ia_bus
port 56 nsew signal output
rlabel metal2 s 82726 299200 82782 300000 6 ia_in
port 57 nsew signal input
rlabel metal2 s 57702 299200 57758 300000 6 is_bus
port 58 nsew signal output
rlabel metal2 s 54574 299200 54630 300000 6 is_in
port 59 nsew signal input
rlabel metal2 s 60830 299200 60886 300000 6 is_oe
port 60 nsew signal output
rlabel metal2 s 1490 299200 1546 300000 6 osc_in
port 61 nsew signal input
rlabel metal2 s 20166 299200 20222 300000 6 phi1_in
port 62 nsew signal input
rlabel metal2 s 29550 299200 29606 300000 6 phi1_out
port 63 nsew signal output
rlabel metal2 s 26422 299200 26478 300000 6 phi2_in
port 64 nsew signal input
rlabel metal2 s 23294 299200 23350 300000 6 phi2_out
port 65 nsew signal output
rlabel metal3 s 0 10752 800 10872 6 sraddr_mux[0]
port 66 nsew signal output
rlabel metal3 s 0 18096 800 18216 6 sraddr_mux[1]
port 67 nsew signal output
rlabel metal3 s 0 25440 800 25560 6 sraddr_mux[2]
port 68 nsew signal output
rlabel metal3 s 0 32784 800 32904 6 sraddr_mux[3]
port 69 nsew signal output
rlabel metal3 s 0 40128 800 40248 6 sraddr_mux[4]
port 70 nsew signal output
rlabel metal3 s 0 47336 800 47456 6 sraddr_mux[5]
port 71 nsew signal output
rlabel metal3 s 0 54680 800 54800 6 sraddr_mux[6]
port 72 nsew signal output
rlabel metal3 s 0 62024 800 62144 6 sraddr_mux[7]
port 73 nsew signal output
rlabel metal3 s 0 3544 800 3664 6 sram_clk1
port 74 nsew signal output
rlabel metal3 s 0 69368 800 69488 6 srdata[0]
port 75 nsew signal input
rlabel metal3 s 0 142536 800 142656 6 srdata[10]
port 76 nsew signal input
rlabel metal3 s 0 149880 800 150000 6 srdata[11]
port 77 nsew signal input
rlabel metal3 s 0 157088 800 157208 6 srdata[12]
port 78 nsew signal input
rlabel metal3 s 0 164432 800 164552 6 srdata[13]
port 79 nsew signal input
rlabel metal3 s 0 171776 800 171896 6 srdata[14]
port 80 nsew signal input
rlabel metal3 s 0 179120 800 179240 6 srdata[15]
port 81 nsew signal input
rlabel metal3 s 0 186464 800 186584 6 srdata[16]
port 82 nsew signal input
rlabel metal3 s 0 193672 800 193792 6 srdata[17]
port 83 nsew signal input
rlabel metal3 s 0 201016 800 201136 6 srdata[18]
port 84 nsew signal input
rlabel metal3 s 0 208360 800 208480 6 srdata[19]
port 85 nsew signal input
rlabel metal3 s 0 76712 800 76832 6 srdata[1]
port 86 nsew signal input
rlabel metal3 s 0 215704 800 215824 6 srdata[20]
port 87 nsew signal input
rlabel metal3 s 0 223048 800 223168 6 srdata[21]
port 88 nsew signal input
rlabel metal3 s 0 230256 800 230376 6 srdata[22]
port 89 nsew signal input
rlabel metal3 s 0 237600 800 237720 6 srdata[23]
port 90 nsew signal input
rlabel metal3 s 0 244944 800 245064 6 srdata[24]
port 91 nsew signal input
rlabel metal3 s 0 252288 800 252408 6 srdata[25]
port 92 nsew signal input
rlabel metal3 s 0 259632 800 259752 6 srdata[26]
port 93 nsew signal input
rlabel metal3 s 0 266840 800 266960 6 srdata[27]
port 94 nsew signal input
rlabel metal3 s 0 274184 800 274304 6 srdata[28]
port 95 nsew signal input
rlabel metal3 s 0 281528 800 281648 6 srdata[29]
port 96 nsew signal input
rlabel metal3 s 0 83920 800 84040 6 srdata[2]
port 97 nsew signal input
rlabel metal3 s 0 288872 800 288992 6 srdata[30]
port 98 nsew signal input
rlabel metal3 s 0 296216 800 296336 6 srdata[31]
port 99 nsew signal input
rlabel metal3 s 0 91264 800 91384 6 srdata[3]
port 100 nsew signal input
rlabel metal3 s 0 98608 800 98728 6 srdata[4]
port 101 nsew signal input
rlabel metal3 s 0 105952 800 106072 6 srdata[5]
port 102 nsew signal input
rlabel metal3 s 0 113296 800 113416 6 srdata[6]
port 103 nsew signal input
rlabel metal3 s 0 120504 800 120624 6 srdata[7]
port 104 nsew signal input
rlabel metal3 s 0 127848 800 127968 6 srdata[8]
port 105 nsew signal input
rlabel metal3 s 0 135192 800 135312 6 srdata[9]
port 106 nsew signal input
rlabel metal2 s 95238 299200 95294 300000 6 sync_bus
port 107 nsew signal output
rlabel metal2 s 98366 299200 98422 300000 6 sync_in
port 108 nsew signal input
rlabel metal4 s 4208 2128 4528 297616 6 vccd1
port 109 nsew power input
rlabel metal4 s 34928 2128 35248 297616 6 vccd1
port 109 nsew power input
rlabel metal4 s 65648 2128 65968 297616 6 vccd1
port 109 nsew power input
rlabel metal4 s 96368 2128 96688 297616 6 vccd1
port 109 nsew power input
rlabel metal4 s 19568 2128 19888 297616 6 vssd1
port 110 nsew ground input
rlabel metal4 s 50288 2128 50608 297616 6 vssd1
port 110 nsew ground input
rlabel metal4 s 81008 2128 81328 297616 6 vssd1
port 110 nsew ground input
rlabel metal2 s 67086 299200 67142 300000 6 ws_bus
port 111 nsew signal output
rlabel metal2 s 63958 299200 64014 300000 6 ws_in
port 112 nsew signal input
rlabel metal2 s 70214 299200 70270 300000 6 ws_oe
port 113 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 100000 300000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 16613596
string GDS_FILE /home/andylithia/openmpw/MPWTRIAL/openlane/hp35_core/runs/hp35_core/results/finishing/hp35_core.magic.gds
string GDS_START 1402616
<< end >>

