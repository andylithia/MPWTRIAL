magic
tech sky130A
magscale 1 2
timestamp 1654559687
<< obsli1 >>
rect 1104 2159 58880 77809
<< obsm1 >>
rect 934 1912 58958 77920
<< metal2 >>
rect 1214 79200 1270 80000
rect 3606 79200 3662 80000
rect 5998 79200 6054 80000
rect 8390 79200 8446 80000
rect 10782 79200 10838 80000
rect 13174 79200 13230 80000
rect 15566 79200 15622 80000
rect 17958 79200 18014 80000
rect 20350 79200 20406 80000
rect 22742 79200 22798 80000
rect 25134 79200 25190 80000
rect 27526 79200 27582 80000
rect 29918 79200 29974 80000
rect 32402 79200 32458 80000
rect 34794 79200 34850 80000
rect 37186 79200 37242 80000
rect 39578 79200 39634 80000
rect 41970 79200 42026 80000
rect 44362 79200 44418 80000
rect 46754 79200 46810 80000
rect 49146 79200 49202 80000
rect 51538 79200 51594 80000
rect 53930 79200 53986 80000
rect 56322 79200 56378 80000
rect 58714 79200 58770 80000
rect 938 0 994 800
rect 2870 0 2926 800
rect 4894 0 4950 800
rect 6918 0 6974 800
rect 8850 0 8906 800
rect 10874 0 10930 800
rect 12898 0 12954 800
rect 14922 0 14978 800
rect 16854 0 16910 800
rect 18878 0 18934 800
rect 20902 0 20958 800
rect 22926 0 22982 800
rect 24858 0 24914 800
rect 26882 0 26938 800
rect 28906 0 28962 800
rect 30930 0 30986 800
rect 32862 0 32918 800
rect 34886 0 34942 800
rect 36910 0 36966 800
rect 38842 0 38898 800
rect 40866 0 40922 800
rect 42890 0 42946 800
rect 44914 0 44970 800
rect 46846 0 46902 800
rect 48870 0 48926 800
rect 50894 0 50950 800
rect 52918 0 52974 800
rect 54850 0 54906 800
rect 56874 0 56930 800
rect 58898 0 58954 800
<< obsm2 >>
rect 940 79144 1158 79200
rect 1326 79144 3550 79200
rect 3718 79144 5942 79200
rect 6110 79144 8334 79200
rect 8502 79144 10726 79200
rect 10894 79144 13118 79200
rect 13286 79144 15510 79200
rect 15678 79144 17902 79200
rect 18070 79144 20294 79200
rect 20462 79144 22686 79200
rect 22854 79144 25078 79200
rect 25246 79144 27470 79200
rect 27638 79144 29862 79200
rect 30030 79144 32346 79200
rect 32514 79144 34738 79200
rect 34906 79144 37130 79200
rect 37298 79144 39522 79200
rect 39690 79144 41914 79200
rect 42082 79144 44306 79200
rect 44474 79144 46698 79200
rect 46866 79144 49090 79200
rect 49258 79144 51482 79200
rect 51650 79144 53874 79200
rect 54042 79144 56266 79200
rect 56434 79144 58658 79200
rect 58826 79144 58952 79200
rect 940 856 58952 79144
rect 1050 734 2814 856
rect 2982 734 4838 856
rect 5006 734 6862 856
rect 7030 734 8794 856
rect 8962 734 10818 856
rect 10986 734 12842 856
rect 13010 734 14866 856
rect 15034 734 16798 856
rect 16966 734 18822 856
rect 18990 734 20846 856
rect 21014 734 22870 856
rect 23038 734 24802 856
rect 24970 734 26826 856
rect 26994 734 28850 856
rect 29018 734 30874 856
rect 31042 734 32806 856
rect 32974 734 34830 856
rect 34998 734 36854 856
rect 37022 734 38786 856
rect 38954 734 40810 856
rect 40978 734 42834 856
rect 43002 734 44858 856
rect 45026 734 46790 856
rect 46958 734 48814 856
rect 48982 734 50838 856
rect 51006 734 52862 856
rect 53030 734 54794 856
rect 54962 734 56818 856
rect 56986 734 58842 856
<< metal3 >>
rect 0 78752 800 78872
rect 59200 78616 60000 78736
rect 0 76712 800 76832
rect 59200 76168 60000 76288
rect 0 74536 800 74656
rect 59200 73720 60000 73840
rect 0 72496 800 72616
rect 59200 71272 60000 71392
rect 0 70320 800 70440
rect 59200 68824 60000 68944
rect 0 68280 800 68400
rect 59200 66512 60000 66632
rect 0 66104 800 66224
rect 0 64064 800 64184
rect 59200 64064 60000 64184
rect 0 61888 800 62008
rect 59200 61616 60000 61736
rect 0 59848 800 59968
rect 59200 59168 60000 59288
rect 0 57672 800 57792
rect 59200 56720 60000 56840
rect 0 55632 800 55752
rect 59200 54408 60000 54528
rect 0 53456 800 53576
rect 59200 51960 60000 52080
rect 0 51416 800 51536
rect 59200 49512 60000 49632
rect 0 49240 800 49360
rect 0 47200 800 47320
rect 59200 47064 60000 47184
rect 0 45024 800 45144
rect 59200 44616 60000 44736
rect 0 42984 800 43104
rect 59200 42168 60000 42288
rect 0 40944 800 41064
rect 59200 39856 60000 39976
rect 0 38768 800 38888
rect 59200 37408 60000 37528
rect 0 36728 800 36848
rect 59200 34960 60000 35080
rect 0 34552 800 34672
rect 0 32512 800 32632
rect 59200 32512 60000 32632
rect 0 30336 800 30456
rect 59200 30064 60000 30184
rect 0 28296 800 28416
rect 59200 27752 60000 27872
rect 0 26120 800 26240
rect 59200 25304 60000 25424
rect 0 24080 800 24200
rect 59200 22856 60000 22976
rect 0 21904 800 22024
rect 59200 20408 60000 20528
rect 0 19864 800 19984
rect 59200 17960 60000 18080
rect 0 17688 800 17808
rect 0 15648 800 15768
rect 59200 15512 60000 15632
rect 0 13472 800 13592
rect 59200 13200 60000 13320
rect 0 11432 800 11552
rect 59200 10752 60000 10872
rect 0 9256 800 9376
rect 59200 8304 60000 8424
rect 0 7216 800 7336
rect 59200 5856 60000 5976
rect 0 5040 800 5160
rect 59200 3408 60000 3528
rect 0 3000 800 3120
rect 0 960 800 1080
rect 59200 1096 60000 1216
<< obsm3 >>
rect 880 78816 59200 78845
rect 880 78672 59120 78816
rect 800 78536 59120 78672
rect 800 76912 59200 78536
rect 880 76632 59200 76912
rect 800 76368 59200 76632
rect 800 76088 59120 76368
rect 800 74736 59200 76088
rect 880 74456 59200 74736
rect 800 73920 59200 74456
rect 800 73640 59120 73920
rect 800 72696 59200 73640
rect 880 72416 59200 72696
rect 800 71472 59200 72416
rect 800 71192 59120 71472
rect 800 70520 59200 71192
rect 880 70240 59200 70520
rect 800 69024 59200 70240
rect 800 68744 59120 69024
rect 800 68480 59200 68744
rect 880 68200 59200 68480
rect 800 66712 59200 68200
rect 800 66432 59120 66712
rect 800 66304 59200 66432
rect 880 66024 59200 66304
rect 800 64264 59200 66024
rect 880 63984 59120 64264
rect 800 62088 59200 63984
rect 880 61816 59200 62088
rect 880 61808 59120 61816
rect 800 61536 59120 61808
rect 800 60048 59200 61536
rect 880 59768 59200 60048
rect 800 59368 59200 59768
rect 800 59088 59120 59368
rect 800 57872 59200 59088
rect 880 57592 59200 57872
rect 800 56920 59200 57592
rect 800 56640 59120 56920
rect 800 55832 59200 56640
rect 880 55552 59200 55832
rect 800 54608 59200 55552
rect 800 54328 59120 54608
rect 800 53656 59200 54328
rect 880 53376 59200 53656
rect 800 52160 59200 53376
rect 800 51880 59120 52160
rect 800 51616 59200 51880
rect 880 51336 59200 51616
rect 800 49712 59200 51336
rect 800 49440 59120 49712
rect 880 49432 59120 49440
rect 880 49160 59200 49432
rect 800 47400 59200 49160
rect 880 47264 59200 47400
rect 880 47120 59120 47264
rect 800 46984 59120 47120
rect 800 45224 59200 46984
rect 880 44944 59200 45224
rect 800 44816 59200 44944
rect 800 44536 59120 44816
rect 800 43184 59200 44536
rect 880 42904 59200 43184
rect 800 42368 59200 42904
rect 800 42088 59120 42368
rect 800 41144 59200 42088
rect 880 40864 59200 41144
rect 800 40056 59200 40864
rect 800 39776 59120 40056
rect 800 38968 59200 39776
rect 880 38688 59200 38968
rect 800 37608 59200 38688
rect 800 37328 59120 37608
rect 800 36928 59200 37328
rect 880 36648 59200 36928
rect 800 35160 59200 36648
rect 800 34880 59120 35160
rect 800 34752 59200 34880
rect 880 34472 59200 34752
rect 800 32712 59200 34472
rect 880 32432 59120 32712
rect 800 30536 59200 32432
rect 880 30264 59200 30536
rect 880 30256 59120 30264
rect 800 29984 59120 30256
rect 800 28496 59200 29984
rect 880 28216 59200 28496
rect 800 27952 59200 28216
rect 800 27672 59120 27952
rect 800 26320 59200 27672
rect 880 26040 59200 26320
rect 800 25504 59200 26040
rect 800 25224 59120 25504
rect 800 24280 59200 25224
rect 880 24000 59200 24280
rect 800 23056 59200 24000
rect 800 22776 59120 23056
rect 800 22104 59200 22776
rect 880 21824 59200 22104
rect 800 20608 59200 21824
rect 800 20328 59120 20608
rect 800 20064 59200 20328
rect 880 19784 59200 20064
rect 800 18160 59200 19784
rect 800 17888 59120 18160
rect 880 17880 59120 17888
rect 880 17608 59200 17880
rect 800 15848 59200 17608
rect 880 15712 59200 15848
rect 880 15568 59120 15712
rect 800 15432 59120 15568
rect 800 13672 59200 15432
rect 880 13400 59200 13672
rect 880 13392 59120 13400
rect 800 13120 59120 13392
rect 800 11632 59200 13120
rect 880 11352 59200 11632
rect 800 10952 59200 11352
rect 800 10672 59120 10952
rect 800 9456 59200 10672
rect 880 9176 59200 9456
rect 800 8504 59200 9176
rect 800 8224 59120 8504
rect 800 7416 59200 8224
rect 880 7136 59200 7416
rect 800 6056 59200 7136
rect 800 5776 59120 6056
rect 800 5240 59200 5776
rect 880 4960 59200 5240
rect 800 3608 59200 4960
rect 800 3328 59120 3608
rect 800 3200 59200 3328
rect 880 2920 59200 3200
rect 800 1296 59200 2920
rect 800 1160 59120 1296
rect 880 1016 59120 1160
rect 880 987 59200 1016
<< metal4 >>
rect 4208 2128 4528 77840
rect 19568 2128 19888 77840
rect 34928 2128 35248 77840
rect 50288 2128 50608 77840
<< obsm4 >>
rect 2635 2347 4128 77349
rect 4608 2347 19488 77349
rect 19968 2347 34848 77349
rect 35328 2347 50208 77349
rect 50688 2347 51461 77349
<< labels >>
rlabel metal2 s 3606 79200 3662 80000 6 COL[0]
port 1 nsew signal input
rlabel metal2 s 5998 79200 6054 80000 6 COL[1]
port 2 nsew signal input
rlabel metal2 s 8390 79200 8446 80000 6 COL[2]
port 3 nsew signal input
rlabel metal2 s 10782 79200 10838 80000 6 COL[3]
port 4 nsew signal input
rlabel metal2 s 13174 79200 13230 80000 6 COL[4]
port 5 nsew signal input
rlabel metal3 s 59200 68824 60000 68944 6 DD[0]
port 6 nsew signal output
rlabel metal3 s 59200 71272 60000 71392 6 DD[1]
port 7 nsew signal output
rlabel metal3 s 59200 73720 60000 73840 6 DD[2]
port 8 nsew signal output
rlabel metal3 s 59200 76168 60000 76288 6 DD[3]
port 9 nsew signal output
rlabel metal3 s 59200 78616 60000 78736 6 DD[4]
port 10 nsew signal output
rlabel metal2 s 1214 79200 1270 80000 6 PWO
port 11 nsew signal input
rlabel metal2 s 15566 79200 15622 80000 6 START
port 12 nsew signal output
rlabel metal2 s 34794 79200 34850 80000 6 bcd_bus
port 13 nsew signal output
rlabel metal2 s 32402 79200 32458 80000 6 bcd_in
port 14 nsew signal input
rlabel metal2 s 37186 79200 37242 80000 6 bcd_oen
port 15 nsew signal output
rlabel metal2 s 46754 79200 46810 80000 6 carry_bus
port 16 nsew signal output
rlabel metal2 s 49146 79200 49202 80000 6 carry_in
port 17 nsew signal input
rlabel metal2 s 51538 79200 51594 80000 6 carry_oen
port 18 nsew signal output
rlabel metal3 s 59200 15512 60000 15632 6 cdiv_rst
port 19 nsew signal input
rlabel metal3 s 59200 51960 60000 52080 6 dbg_arc_a1
port 20 nsew signal output
rlabel metal3 s 59200 54408 60000 54528 6 dbg_arc_b1
port 21 nsew signal output
rlabel metal3 s 59200 44616 60000 44736 6 dbg_arc_dummy
port 22 nsew signal input
rlabel metal3 s 59200 47064 60000 47184 6 dbg_arc_t1
port 23 nsew signal output
rlabel metal3 s 59200 49512 60000 49632 6 dbg_arc_t4
port 24 nsew signal output
rlabel metal3 s 59200 27752 60000 27872 6 dbg_ctc_kdn
port 25 nsew signal output
rlabel metal3 s 59200 30064 60000 30184 6 dbg_ctc_q[0]
port 26 nsew signal output
rlabel metal3 s 59200 32512 60000 32632 6 dbg_ctc_q[1]
port 27 nsew signal output
rlabel metal3 s 59200 34960 60000 35080 6 dbg_ctc_q[2]
port 28 nsew signal output
rlabel metal3 s 59200 37408 60000 37528 6 dbg_ctc_q[3]
port 29 nsew signal output
rlabel metal3 s 59200 39856 60000 39976 6 dbg_ctc_q[4]
port 30 nsew signal output
rlabel metal3 s 59200 42168 60000 42288 6 dbg_ctc_q[5]
port 31 nsew signal output
rlabel metal3 s 59200 25304 60000 25424 6 dbg_ctc_state1
port 32 nsew signal output
rlabel metal2 s 42890 0 42946 800 6 dbg_disable_arc
port 33 nsew signal input
rlabel metal2 s 44914 0 44970 800 6 dbg_disable_ctc
port 34 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 dbg_disable_rom
port 35 nsew signal input
rlabel metal3 s 59200 56720 60000 56840 6 dbg_dsbf[0]
port 36 nsew signal output
rlabel metal3 s 59200 59168 60000 59288 6 dbg_dsbf[1]
port 37 nsew signal output
rlabel metal3 s 59200 61616 60000 61736 6 dbg_dsbf[2]
port 38 nsew signal output
rlabel metal3 s 59200 64064 60000 64184 6 dbg_dsbf[3]
port 39 nsew signal output
rlabel metal3 s 59200 66512 60000 66632 6 dbg_dsbf[4]
port 40 nsew signal output
rlabel metal3 s 59200 20408 60000 20528 6 dbg_force_data
port 41 nsew signal input
rlabel metal3 s 59200 17960 60000 18080 6 dbg_internal_cdiv
port 42 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 dbg_rom_roe[0]
port 43 nsew signal output
rlabel metal2 s 38842 0 38898 800 6 dbg_rom_roe[1]
port 44 nsew signal output
rlabel metal2 s 40866 0 40922 800 6 dbg_rom_roe[2]
port 45 nsew signal output
rlabel metal2 s 16854 0 16910 800 6 dbg_romdata[0]
port 46 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 dbg_romdata[1]
port 47 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 dbg_romdata[2]
port 48 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 dbg_romdata[3]
port 49 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 dbg_romdata[4]
port 50 nsew signal input
rlabel metal2 s 26882 0 26938 800 6 dbg_romdata[5]
port 51 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 dbg_romdata[6]
port 52 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 dbg_romdata[7]
port 53 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 dbg_romdata[8]
port 54 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 dbg_romdata[9]
port 55 nsew signal input
rlabel metal3 s 59200 5856 60000 5976 6 dbg_sram_cksel[0]
port 56 nsew signal input
rlabel metal3 s 59200 8304 60000 8424 6 dbg_sram_cksel[1]
port 57 nsew signal input
rlabel metal3 s 59200 10752 60000 10872 6 dbg_sram_cksel[2]
port 58 nsew signal input
rlabel metal3 s 59200 22856 60000 22976 6 dbg_sram_csb1
port 59 nsew signal input
rlabel metal3 s 59200 1096 60000 1216 6 dbg_sram_wrmode[0]
port 60 nsew signal input
rlabel metal3 s 59200 3408 60000 3528 6 dbg_sram_wrmode[1]
port 61 nsew signal input
rlabel metal2 s 41970 79200 42026 80000 6 ia_bus
port 62 nsew signal output
rlabel metal2 s 39578 79200 39634 80000 6 ia_in
port 63 nsew signal input
rlabel metal2 s 44362 79200 44418 80000 6 ia_oen
port 64 nsew signal output
rlabel metal2 s 20350 79200 20406 80000 6 is_bus
port 65 nsew signal output
rlabel metal2 s 17958 79200 18014 80000 6 is_in
port 66 nsew signal input
rlabel metal2 s 22742 79200 22798 80000 6 is_oen
port 67 nsew signal output
rlabel metal2 s 48870 0 48926 800 6 osc_in
port 68 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 phi1_in
port 69 nsew signal input
rlabel metal2 s 56874 0 56930 800 6 phi1_out
port 70 nsew signal output
rlabel metal2 s 54850 0 54906 800 6 phi2_in
port 71 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 phi2_out
port 72 nsew signal output
rlabel metal2 s 58898 0 58954 800 6 phi_oen
port 73 nsew signal output
rlabel metal2 s 938 0 994 800 6 sraddr_in[0]
port 74 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 sraddr_in[1]
port 75 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 sraddr_in[2]
port 76 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 sraddr_in[3]
port 77 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 sraddr_in[4]
port 78 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 sraddr_in[5]
port 79 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 sraddr_in[6]
port 80 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 sraddr_in[7]
port 81 nsew signal input
rlabel metal3 s 0 960 800 1080 6 sraddr_mux[0]
port 82 nsew signal output
rlabel metal3 s 0 3000 800 3120 6 sraddr_mux[1]
port 83 nsew signal output
rlabel metal3 s 0 5040 800 5160 6 sraddr_mux[2]
port 84 nsew signal output
rlabel metal3 s 0 7216 800 7336 6 sraddr_mux[3]
port 85 nsew signal output
rlabel metal3 s 0 9256 800 9376 6 sraddr_mux[4]
port 86 nsew signal output
rlabel metal3 s 0 11432 800 11552 6 sraddr_mux[5]
port 87 nsew signal output
rlabel metal3 s 0 13472 800 13592 6 sraddr_mux[6]
port 88 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 sraddr_mux[7]
port 89 nsew signal output
rlabel metal3 s 59200 13200 60000 13320 6 sram_clk1
port 90 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 srdata[0]
port 91 nsew signal input
rlabel metal3 s 0 38768 800 38888 6 srdata[10]
port 92 nsew signal input
rlabel metal3 s 0 40944 800 41064 6 srdata[11]
port 93 nsew signal input
rlabel metal3 s 0 42984 800 43104 6 srdata[12]
port 94 nsew signal input
rlabel metal3 s 0 45024 800 45144 6 srdata[13]
port 95 nsew signal input
rlabel metal3 s 0 47200 800 47320 6 srdata[14]
port 96 nsew signal input
rlabel metal3 s 0 49240 800 49360 6 srdata[15]
port 97 nsew signal input
rlabel metal3 s 0 51416 800 51536 6 srdata[16]
port 98 nsew signal input
rlabel metal3 s 0 53456 800 53576 6 srdata[17]
port 99 nsew signal input
rlabel metal3 s 0 55632 800 55752 6 srdata[18]
port 100 nsew signal input
rlabel metal3 s 0 57672 800 57792 6 srdata[19]
port 101 nsew signal input
rlabel metal3 s 0 19864 800 19984 6 srdata[1]
port 102 nsew signal input
rlabel metal3 s 0 59848 800 59968 6 srdata[20]
port 103 nsew signal input
rlabel metal3 s 0 61888 800 62008 6 srdata[21]
port 104 nsew signal input
rlabel metal3 s 0 64064 800 64184 6 srdata[22]
port 105 nsew signal input
rlabel metal3 s 0 66104 800 66224 6 srdata[23]
port 106 nsew signal input
rlabel metal3 s 0 68280 800 68400 6 srdata[24]
port 107 nsew signal input
rlabel metal3 s 0 70320 800 70440 6 srdata[25]
port 108 nsew signal input
rlabel metal3 s 0 72496 800 72616 6 srdata[26]
port 109 nsew signal input
rlabel metal3 s 0 74536 800 74656 6 srdata[27]
port 110 nsew signal input
rlabel metal3 s 0 76712 800 76832 6 srdata[28]
port 111 nsew signal input
rlabel metal3 s 0 78752 800 78872 6 srdata[29]
port 112 nsew signal input
rlabel metal3 s 0 21904 800 22024 6 srdata[2]
port 113 nsew signal input
rlabel metal3 s 0 24080 800 24200 6 srdata[3]
port 114 nsew signal input
rlabel metal3 s 0 26120 800 26240 6 srdata[4]
port 115 nsew signal input
rlabel metal3 s 0 28296 800 28416 6 srdata[5]
port 116 nsew signal input
rlabel metal3 s 0 30336 800 30456 6 srdata[6]
port 117 nsew signal input
rlabel metal3 s 0 32512 800 32632 6 srdata[7]
port 118 nsew signal input
rlabel metal3 s 0 34552 800 34672 6 srdata[8]
port 119 nsew signal input
rlabel metal3 s 0 36728 800 36848 6 srdata[9]
port 120 nsew signal input
rlabel metal2 s 53930 79200 53986 80000 6 sync_bus
port 121 nsew signal output
rlabel metal2 s 56322 79200 56378 80000 6 sync_in
port 122 nsew signal input
rlabel metal2 s 58714 79200 58770 80000 6 sync_oen
port 123 nsew signal output
rlabel metal4 s 4208 2128 4528 77840 6 vccd1
port 124 nsew power input
rlabel metal4 s 34928 2128 35248 77840 6 vccd1
port 124 nsew power input
rlabel metal4 s 19568 2128 19888 77840 6 vssd1
port 125 nsew ground input
rlabel metal4 s 50288 2128 50608 77840 6 vssd1
port 125 nsew ground input
rlabel metal2 s 27526 79200 27582 80000 6 ws_bus
port 126 nsew signal output
rlabel metal2 s 25134 79200 25190 80000 6 ws_in
port 127 nsew signal input
rlabel metal2 s 29918 79200 29974 80000 6 ws_oen
port 128 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 60000 80000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9240214
string GDS_FILE /home/andylithia/openmpw/MPWTRIAL/openlane/hp35_core/runs/hp35_core/results/finishing/hp35_core.magic.gds
string GDS_START 1173226
<< end >>

