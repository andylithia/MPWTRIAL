module rom_tb;




endmodule